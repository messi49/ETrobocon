/*
 *   TOPPERS Software
 *       Toyohashi Open Platform for Embedded Real-Time Systems
 *  
 *   Copyright (C) 2010-2012 by Embedded and Real-Time Systems Laboratory
 *               Graduate School of Information Science, Nagoya Univ., JAPAN
 *  
 *   �嵭����Ԥϡ��ʲ���(1)��(4)�ξ������������˸¤ꡤ�ܥ��եȥ���
 *   �����ܥ��եȥ���������Ѥ�����Τ�ޤࡥ�ʲ�Ʊ���ˤ���ѡ�ʣ������
 *   �ѡ������ۡʰʲ������ѤȸƤ֡ˤ��뤳�Ȥ�̵���ǵ������롥
 *   (1) �ܥ��եȥ������򥽡��������ɤη������Ѥ�����ˤϡ��嵭������
 *       ��ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ��꤬�����Τޤޤη��ǥ���
 *       ����������˴ޤޤ�Ƥ��뤳�ȡ�
 *   (2) �ܥ��եȥ������򡤥饤�֥������ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ�����Ǻ����ۤ�����ˤϡ������ۤ�ȼ���ɥ�����ȡ�����
 *       �ԥޥ˥奢��ʤɡˤˡ��嵭�����ɽ�����������Ѿ�浪��Ӳ���
 *       ��̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *   (3) �ܥ��եȥ������򡤵�����Ȥ߹���ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ��ʤ����Ǻ����ۤ�����ˤϡ����Τ����줫�ξ�����������
 *       �ȡ�
 *     (a) �����ۤ�ȼ���ɥ�����ȡ����Ѽԥޥ˥奢��ʤɡˤˡ��嵭����
 *         �ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *     (b) �����ۤη��֤��̤�������ˡ�ˤ�äơ�TOPPERS�ץ������Ȥ�
 *         ��𤹤뤳�ȡ�
 *   (4) �ܥ��եȥ����������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������뤤���ʤ�»
 *       ������⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ����դ��뤳�ȡ�
 *       �ޤ����ܥ��եȥ������Υ桼���ޤ��ϥ���ɥ桼������Τ����ʤ���
 *       ͳ�˴�Ť����ᤫ��⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ�
 *       ���դ��뤳�ȡ�
 *  
 *   �ܥ��եȥ������ϡ�̵�ݾڤ��󶡤���Ƥ����ΤǤ��롥�嵭����Ԥ�
 *   ���TOPPERS�ץ������Ȥϡ��ܥ��եȥ������˴ؤ��ơ�����λ�����Ū
 *   ���Ф���Ŭ������ޤ�ơ������ʤ��ݾڤ�Ԥ�ʤ����ޤ����ܥ��եȥ���
 *   �������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������������ʤ�»���˴ؤ��Ƥ⡤��
 *   ����Ǥ�����ʤ���
 *
 */

/*
 *  ����ץ�ץ��������
 */


/*
 *  fujiya
 *	�ǥ����ץ쥤ɽ����
 */

signature sPrintDisplayControl{
 
    //structure��
    void print_str(void);

    //kp,ki,kd
    void print_k([in]const char* string1, [in] int16_t value1);
	

    //�ͤ���
    void print1([in] int16_t value1);
    void print2([in] int16_t value1, [in] int16_t value2);
    void print3([in] int16_t value1, [in] int16_t value2, [in] int16_t value3);
    void print4([in] int16_t value1, [in] int16_t value2, [in] int16_t value3, [in] int16_t value4);
    void print5([in] int16_t value1,[in] int16_t value2,[in] int16_t value3,[in] int16_t value4,[in] int16_t value5);

    void print6([in] int16_t value1,[in] int16_t value2,[in] int16_t value3,[in] int16_t value4,[in] int16_t value5, [in]int16_t value6);
    void print7([in] int16_t value1,[in] int16_t value2,[in] int16_t value3,[in] int16_t value4,[in] int16_t value5, [in]int16_t value6, [in]int16_t value7);



    //�ͤ�String
    void printS1([in]const char* string1, [in] int16_t value1);
    void printS2([in]const char* string1, [in] int16_t value1,[in]const char* string2, [in] int16_t value2);
    void printS3([in]const char* string1, [in] int16_t value1, [in]const char* string2, [in] int16_t value2, [in]const char* string3, [in] int16_t value3);
};

[singleton]
celltype tPrintDisplayTaskBody{
	entry sPrintDisplayControl ePrintDisplayControl; // �������ѥ�᡼�����åȤμ�����

	call sDisplay cDisplay;
};
/*
 *  PID���楿���� by no- (2013/08/18)
 */
signature sPIDControl{
  void getPIDValue( [in]uint16_t light, [in] uint16_t VAR_lightThreshold,[out] float32_t *turn_f);
  void getKValue([out] float32_t *kp, [out]float32_t *ki, [out]float32_t *kd);
  void setKValue([in] uint8_t kind, [in] float32_t value);
};

[singleton]
celltype tPIDControllerTaskBody{
   require tKernel.eKernel;
   entry sPIDControl ePIDControl;

  var{
    float32_t kp=0.6;
    float32_t ki=0;
    float32_t kd=0.2;

    float32_t integral=0;
    float32_t diff0=0;
    float32_t diff1=0;
    float32_t DELTAT=0.010;  //0.004?
  };

};

/*
 *  �������楿����
 */
/*
 *  �����������åȳ�����
 */
signature sTailController{
    void setAngle([in] int32_t angle);
    void getAngle([out] int32_t *angle);
	//void setStopAngle([in] int32_t angle);
	//void getStopAngle([out] int32_t *angle);
	//void setDriveAngle([in] int32_t angle);
	//void getDriveAngle([out] int32_t *angle);
	void signalStop(void);
	void signalStart(void);
    void calibrate(void);
};

[singleton]
celltype tTailControllerTaskBody{
	require tKernel.eKernel;
	
	entry sTaskBody eBody;        // ���������Τμ�����
	entry sTailController eTailController; // �����������åȳ�����μ�����
	
	call sMotor cTailMotor;       // �����⡼���θƤӸ�
	
	attr{
		int32_t tailAngleStop;
		int32_t tailAngleDrive;
		float32_t kp;
		int8_t maxPwm;
		int8_t minPwm;
	};
	var{
		int32_t targetAngle;
		
	};
};

/*
 *  �Х�󥵥�����
 */
/*
 *  �Х�󥵥������ѥ�᡼�����åȤΥ����˥���
 */
signature sBalancerControl{
	void setSpeed([in] int16_t speed);
	void getSpeed([out] int16_t *speed);
	void setTurn([in] int16_t turn);
	void getTurn([out] int16_t *turn);
        void calibrate(void);
};

[singleton]
celltype tBalancerTaskBody{
	require tKernel.eKernel;
	
	entry sTaskBody eBody;     // ���������Τμ�����
	entry sBalancerControl eBalancerControl; // �Х�󥵥������ѥ�᡼�����åȤμ�����
	call sMotor cRightMotor;  // ���⡼���θƤӸ�
	call sMotor cLeftMotor;   // ���⡼���θƤӸ�
	call sSensor cGyroSensor; // ���㥤���󥵤θƤӸ�
	call sBattery cBattery;   // �Хåƥꥻ�󥵤θƤӸ�
	call sBalancer cBalancer; // �Х�󥵤θƤӸ�

	//fujiya �ǥХå��ѡ��ǥ����ץ쥤ɽ��
	call sPrintDisplayControl cPrintDisplayControl; 
	
	attr{
		int16_t maxSpeed;
		int16_t minSpeed;
	};
	var{
		uint16_t gyroOffset;
		int16_t speed;
		int16_t turn;
        	int32_t count = 0;

	};
};

/*
 *  �饤��ȥ졼��������
 */
/*
 *  �饤��ȥ졼���������ѥ�᡼�����åȤΥ����˥���
 */
signature sLinetracerControl{
    void setLightThreshold ([in] uint8_t color, [in] uint16_t light);
    void getLightThreshold ([in] uint8_t color, [out] uint16_t *light);
    void setEdge([in] int8_t edge);
    void getEdge([out] int8_t *edge);


};

[singleton]
celltype tLinetracerTaskBody{
	require tKernel.eKernel;

	entry sTaskBody eBody;     // ���������Τμ�����
	entry sLinetracerControl eLinetracerControl; // �������ѥ�᡼�����åȤμ�����
	call sSensor cLightSensor; // �����󥵤θƤӸ�
	call sSensorControl cLightSensorControl; // ����������θƤӸ�
	call sBalancerControl cBalancerControl; // �Х�󥵥������ѥ�᡼�����åȤθƤӸ�

	call sPIDControl cPIDControl; //no(2013/08/18)
	
	//fujiya���ǥХå��ѡ��ǥ����ץ쥤ɽ��
	call sPrintDisplayControl cPrintDisplayControl; 
	call sMotor cRightMotor; // �⡼���β�ž���μ����Τ���(2011/08/17 itwu added)
  	call sMotor cLeftMotor; // �⡼���β�ž���μ����Τ���(2011/08/17 itwu added)

	call sCyclic cBalancerTask;     // �Х�󥵥������θƤӸ�
	call sCyclic cLinetracerTask;    // �饤��ȥ졼���������θƤӸ�


	attr{
		int16_t maxTurn;
		int16_t minTurn;
      
	};

	var{
		uint16_t lightThreshold;
      	int8_t  edge;
        uint16_t black;
        uint16_t white;
        int32_t count = 0;

        float32_t xx=0;
        float32_t yy =0;
        float32_t sita=0;
        int32_t preLeft = 0;
        int32_t preRight = 0;
	};
};
	
/*
 *  added by no
 *	�ܥ��������
 */

signature sButtonSetValue{
 
    //�ͤ���
    void kvalue(void);
    void threshold(void);
    void speed(void);
    void tailAngle(void);
  
};

[singleton]
celltype tButtonSetTaskBody{
	require tKernel.eKernel;
	entry sButtonSetValue eButtonSetValue; // �������ѥ�᡼�����åȤμ�����

	call sButton cButton;
	call sDisplay cDisplay;
	call sPIDControl cPIDControl; /*added by no 13.08.26*/
	call sLinetracerControl cLinetracerControl; /*added by no 13.08.27*/
	call sBalancerControl cBalancerControl; /*added by no*/
	call sTailController cTailController;
	call sPrintDisplayControl cPrintDisplayControl; 
	call sSensor cTouchSensor;
};

/*
 *  messi
 *	�����ϥ�����
 */

signature sGetLogControl{
	void portOpen(void); 
};

 [singleton]
celltype tGetLogTaskBody{
	require tKernel.eKernel;
	
	entry sTaskBody eBody;     // ���������Τμ�����
	entry sGetLogControl eGetLogControl; // �������ѥ�᡼�����åȤμ�����

	call sSerialPort cSerialPort; // ���ꥢ��ݡ��ȤθƤӸ�
    call sSysLog cSysLog;
	call sLinetracerControl cLinetracerControl;
    call sBalancerControl cBalancerControl;
    call sTailController cTailController;
    call sSemaphore cSemaphore; // ���ޥե��θƤӸ�

    //messi added
	call sSensor cLightSensor; // �����󥵤θƤӸ�

	//fujiy added
	call sMotor cRightMotor; // �⡼���β�ž���μ����Τ���
  	call sMotor cLeftMotor; // �⡼���β�ž���μ����Τ���


};




/*
 *  ��������������
 */
[singleton]
celltype tStarterTaskBody{
	require tKernel.eKernel;  // �����ͥ�Υ����ӥ�������
	
	entry sTaskBody eBody;        // ���������Τμ�����

	call sCyclic cTailControllerTask;     // �������楿�����θƤӸ�
	call sCyclic cBalancerTask;     // �Х�󥵥������θƤӸ�
	call sCyclic cLinetracerTask;    // �饤��ȥ졼���������θƤӸ�
	call sCyclic cGetLogTask;		//Log���ϥ�����
	call sTailController cTailController; // �����������åȳ�����θƤӸ�

	call sSemaphore cSemaphore; // ���ޥե��θƤӸ�
	//[optional] call sSensor cTouchSensor;
	
	// fujiya:���ǥХå���
	call sPrintDisplayControl cPrintDisplayControl; 

	// added by no �ܥ���������
	call sButtonSetValue cButtonSetValue;
	call sBattery cBattery;   // �Хåƥꥻ�󥵤θƤӸ�
	call sSensor cLightSensor;
	call sSensor cTouchSensor;
	call sBalancerControl cBalancerControl; // �Х�󥵥������ѥ�᡼�����åȤθƤӸ�
	call sLinetracerControl cLinetracerControl;

	call sGetLogControl cGetLogControl;
};


/*
 *  ���ޥ�ɼ���������
 */
[singleton]
celltype tGetCommandTaskBody{
	require tKernel.eKernel;
	
	entry sTaskBody eBody;     // ���������Τμ�����

	call sSerialPort cSerialPort; // ���ꥢ��ݡ��ȤθƤӸ�
    call sSysLog cSysLog;
	call sLinetracerControl cLinetracerControl;
    call sBalancerControl cBalancerControl;
    call sTailController cTailController;
    call sSemaphore cSemaphore; // ���ޥե��θƤӸ�
	

    //fujiya
	call sSensor cTouchSensor;
	call sPrintDisplayControl cPrintDisplayControl; 
	call sCyclic cBalancerTask;     // �Х�󥵥������θƤӸ�
	call sCyclic cLinetracerTask;    // �饤��ȥ졼���������θƤӸ�

	var{
        int32_t parameter = 0;
        int8_t  sign = 1;
	};
};



/*
 *   TOPPERS Software
 *       Toyohashi Open Platform for Embedded Real-Time Systems
 *  
 *   Copyright (C) 2010-2012 by Embedded and Real-Time Systems Laboratory
 *               Graduate School of Information Science, Nagoya Univ., JAPAN
 *  
 *   �嵭����Ԥϡ��ʲ���(1)��(4)�ξ������������˸¤ꡤ�ܥ��եȥ���
 *   �����ܥ��եȥ���������Ѥ�����Τ�ޤࡥ�ʲ�Ʊ���ˤ���ѡ�ʣ������
 *   �ѡ������ۡʰʲ������ѤȸƤ֡ˤ��뤳�Ȥ�̵���ǵ������롥
 *   (1) �ܥ��եȥ������򥽡��������ɤη������Ѥ�����ˤϡ��嵭������
 *       ��ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ��꤬�����Τޤޤη��ǥ���
 *       ����������˴ޤޤ�Ƥ��뤳�ȡ�
 *   (2) �ܥ��եȥ������򡤥饤�֥������ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ�����Ǻ����ۤ�����ˤϡ������ۤ�ȼ���ɥ�����ȡ�����
 *       �ԥޥ˥奢��ʤɡˤˡ��嵭�����ɽ�����������Ѿ�浪��Ӳ���
 *       ��̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *   (3) �ܥ��եȥ������򡤵�����Ȥ߹���ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ��ʤ����Ǻ����ۤ�����ˤϡ����Τ����줫�ξ�����������
 *       �ȡ�
 *     (a) �����ۤ�ȼ���ɥ�����ȡ����Ѽԥޥ˥奢��ʤɡˤˡ��嵭����
 *         �ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *     (b) �����ۤη��֤��̤�������ˡ�ˤ�äơ�TOPPERS�ץ������Ȥ�
 *         ��𤹤뤳�ȡ�
 *   (4) �ܥ��եȥ����������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������뤤���ʤ�»
 *       ������⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ����դ��뤳�ȡ�
 *       �ޤ����ܥ��եȥ������Υ桼���ޤ��ϥ���ɥ桼������Τ����ʤ���
 *       ͳ�˴�Ť����ᤫ��⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ�
 *       ���դ��뤳�ȡ�
 *  
 *   �ܥ��եȥ������ϡ�̵�ݾڤ��󶡤���Ƥ����ΤǤ��롥�嵭����Ԥ�
 *   ���TOPPERS�ץ������Ȥϡ��ܥ��եȥ������˴ؤ��ơ�����λ�����Ū
 *   ���Ф���Ŭ������ޤ�ơ������ʤ��ݾڤ�Ԥ�ʤ����ޤ����ܥ��եȥ���
 *   �������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������������ʤ�»���˴ؤ��Ƥ⡤��
 *   ����Ǥ�����ʤ���
 *
 */

/*
 *  �Ȥ߾夲����
 */
/*
 *  �����ƥ������
 */
cell tSerialPort SerialPort1 {
	/* �ƤӸ��η�� */
	cSIOPort = SIOPortTarget.eSIOPort;
	receiveBufferSize = 256;
	sendBufferSize = 256;
};

cell tSysLog SysLog {
	/* �ƤӸ��η�� */
	cPutLog = PutLogTarget.ePutLog;
	logBufferSize = 32;
};

cell tLogTask LogTask {
	/* �ƤӸ��η�� */
	cSerialPort = SerialPort1.eSerialPort;
	cnSerialPort = SerialPort1.enSerialPort;
	cSysLog = SysLog.eSysLog;
	cPutLog = PutLogTarget.ePutLog;
	/* °�������� */
	taskAttribute = C_EXP("TA_ACT");
	priority = 3;
	stackSize = LogTaskStackSize;
	
};

/*
 *  ����
 */
cell tGyroSensor GyroSensor{
	portNumber = NXT_PORT_S1;
	cAvrSensor = AVR.eAvrSensor;
};

cell tSonicSensor SonicSensor{
	portNumber = NXT_PORT_S2;
	cAvrSensor = AVR.eAvrSensor;
};

cell tLightSensor LightSensor{
	portNumber = NXT_PORT_S3;
	cAvrSensor = AVR.eAvrSensor;
};

cell tTouchSensor TouchSensor{
	portNumber = NXT_PORT_S4;
	cAvrSensor = AVR.eAvrSensor;
};

cell tSensorDriver SensorDriver{
	ciSensorDriver[0] = GyroSensor.eiSensorDriver;
	ciSensorDriver[1] = SonicSensor.eiSensorDriver;
	ciSensorDriver[2] = LightSensor.eiSensorDriver;
	ciSensorDriver[3] = TouchSensor.eiSensorDriver;
};

/*
 *  �⡼��
 */
cell tMotor TailMotor{
	portNumber = NXT_PORT_A;
	cAvrMotor = AVR.eAvrMotor;
};

cell tMotor RightMotor{
	portNumber = NXT_PORT_B;
	cAvrMotor = AVR.eAvrMotor;
};

cell tMotor LeftMotor{
	portNumber = NXT_PORT_C;
	cAvrMotor = AVR.eAvrMotor;
};

cell tRotaryEncoder RotaryEncoder{
	ciMotorInterrupt[0] = TailMotor.eiMotorInterrupt;
	ciMotorInterrupt[1] = RightMotor.eiMotorInterrupt;
	ciMotorInterrupt[2] = LeftMotor.eiMotorInterrupt;
};

/*
 *  �Хåƥꥻ��
 */
cell tBattery Battery{
	cAvrBattery = AVR.eAvrBattery;
};

/*
 *  �ǥ����ץ쥤
 */
cell tDisplay Display{
};

/*
 *  �������
 */
cell tSound Sound{
};

/*
 *  �Х�󥵡ʥ饤�֥���
 */
cell tBalancer Balancer{
};

/*
 *  ASP�����ͥ�
 */
cell tKernel ASPKernel{
};

/*
 *  PID���楿���� by no(13/08/18)
 */
cell tPIDControllerTaskBody PIDControllerTaskBody{
	//kp = 0.6;	//0.75, 0.6 , 0.36
	//ki = 0;  	//0, 0.4 , 1.2 (0.00->0.01->0.06)
	//kd = 0.2;	//0.85, 0.2 , 0.027

};

/*
 *  �������楿����
 */
cell tTailControllerTaskBody TailControllerTaskBody{
	cTailMotor = TailMotor.eMotor;       // �����⡼���θƤӸ�
	
	tailAngleStop = 106; //90����Ω
	tailAngleDrive = 60; //60:
	kp = 2.5;
	maxPwm = 60;
	minPwm = -60;
};
cell tCyclicTask TailControllerTask{
	cBody = TailControllerTaskBody.eBody;

	cyclicAttribute = C_EXP("TA_NULL");
	cyclicTime = 4;
	cyclicPhase = 1;
	priority = 5;
	stackSize = 512;
};

/*
 *  �Х�󥵥�����
 */
cell tBalancerTaskBody BalancerTaskBody{
	cRightMotor = RightMotor.eMotor;
	cLeftMotor = LeftMotor.eMotor;
	cGyroSensor = GyroSensor.eSensor;
	cBattery = Battery.eBattery;
	cBalancer = Balancer.eBalancer;
	
	//fujiya
	cPrintDisplayControl = PrintDisplayTaskBody.ePrintDisplayControl;

	maxSpeed = 100;
	minSpeed = -100;

};

cell tCyclicTask BalancerTask{
	cBody = BalancerTaskBody.eBody;

	cyclicAttribute = C_EXP("TA_NULL");
	cyclicTime = 4;
	cyclicPhase = 1;
	priority = 1;
	stackSize = 1024;
};

/*
 *  �饤��ȥ졼��������
 */
cell tLinetracerTaskBody LinetracerTaskBody{
	cLightSensor = LightSensor.eSensor;
	cLightSensorControl = LightSensor.eSensorControl;
	cBalancerControl = BalancerTaskBody.eBalancerControl;

	cPIDControl = PIDControllerTaskBody.ePIDControl; //no(13/08/18)
	//fujiya
	cPrintDisplayControl = PrintDisplayTaskBody.ePrintDisplayControl;

	//fujiya from zukky program
	cRightMotor = RightMotor.eMotor;// �⡼���β�ž���μ����Τ���(2011/08/17 itwu added)
 	cLeftMotor = LeftMotor.eMotor;// �⡼���β�ž���μ����Τ���(2011/08/17 itwu added)

 	cBalancerTask = BalancerTask.eCyclic;
	cLinetracerTask = LinetracerTask.eCyclic;
  
	maxTurn = 100;
	minTurn = -100;

};

cell tCyclicTask LinetracerTask{
	cBody = LinetracerTaskBody.eBody;

	cyclicAttribute = C_EXP("TA_NULL");
	cyclicTime = 10;
	cyclicPhase = 1;
	priority = 4;
	stackSize = 512;
};

/*
 *  �������ȥ����ʥ��ѥ��ޥե�
 */
cell tSemaphore StartSemaphore{
	attribute = C_EXP("TA_NULL");
    	count = 0;  /* ����񸻿���0 */
    	max = 1;    /* ����񸻿���1 */
};

/*
 *  ��������������
 */
cell tStarterTaskBody StarterTaskBody{
    /*
     *  �����������ε�ư
     */
	cTailControllerTask = TailControllerTask.eCyclic;
	cBalancerTask = BalancerTask.eCyclic;
	cLinetracerTask = LinetracerTask.eCyclic;
	cTailController = TailControllerTaskBody.eTailController;
	cGetLogTask = GetLogTask.eCyclic;

    cSemaphore = StartSemaphore.eSemaphore;
	//fujiya
	cPrintDisplayControl = PrintDisplayTaskBody.ePrintDisplayControl;

	//added by no 2013.08.26
	cButtonSetValue = ButtonSetTaskBody.eButtonSetValue;

	cBattery = Battery.eBattery;
	cLightSensor = LightSensor.eSensor;
	cTouchSensor = TouchSensor.eSensor;
	cBalancerControl = BalancerTaskBody.eBalancerControl;
	cLinetracerControl = LinetracerTaskBody.eLinetracerControl;

	cGetLogControl = GetLogTaskBody.eGetLogControl;
};

cell tTask StarterTask{
	cBody = StarterTaskBody.eBody;

	taskAttribute = C_EXP("TA_ACT");
	priority = 6;
	stackSize = 1024;
};

/*
 *  ���ޥ�ɼ���������
 */
cell tGetCommandTaskBody GetCommandTaskBody{
	cSerialPort = SerialPort1.eSerialPort;
        cSysLog = SysLog.eSysLog;
 	cLinetracerControl = LinetracerTaskBody.eLinetracerControl;
        cBalancerControl = BalancerTaskBody.eBalancerControl;
	cTailController = TailControllerTaskBody.eTailController;

    	cSemaphore = StartSemaphore.eSemaphore;


	//fujiya
	cPrintDisplayControl = PrintDisplayTaskBody.ePrintDisplayControl;
        cTouchSensor = TouchSensor.eSensor;

        	cBalancerTask = BalancerTask.eCyclic;
	cLinetracerTask = LinetracerTask.eCyclic;
};

cell tTask GetCommandTask{
	cBody = GetCommandTaskBody.eBody;

	taskAttribute = C_EXP("TA_ACT");
	priority = 5;
	stackSize = 1024;
};

/*
 *  fujiya
 *	�ǥ����ץ쥤ɽ��
 */
cell tPrintDisplayTaskBody PrintDisplayTaskBody {
	cDisplay = Display.eDisplay;
};


/*
 *  �ܥ��������ѥ�����
 */
cell tButtonSetTaskBody ButtonSetTaskBody{
	cButton = Button.eButton;       // �ܥ���θƤӸ�
	cTouchSensor = TouchSensor.eSensor;
	cDisplay = Display.eDisplay;  //Display�θƤӸ�
	cPIDControl = PIDControllerTaskBody.ePIDControl; //no(13/08/26)
	cLinetracerControl = LinetracerTaskBody.eLinetracerControl; //no(13/08/26)
	cBalancerControl = BalancerTaskBody.eBalancerControl; //no
	cTailController = TailControllerTaskBody.eTailController; //no
	cPrintDisplayControl = PrintDisplayTaskBody.ePrintDisplayControl;
	
};

/*
 *  messi
 *  �����ϥ�����
 */
cell tGetLogTaskBody GetLogTaskBody{
	cSerialPort = SerialPort1.eSerialPort;
    cSysLog = SysLog.eSysLog;
	cLinetracerControl = LinetracerTaskBody.eLinetracerControl;
    cBalancerControl = BalancerTaskBody.eBalancerControl;
	cTailController = TailControllerTaskBody.eTailController;

    cSemaphore = StartSemaphore.eSemaphore;

    cLightSensor = LightSensor.eSensor;

    //fujiya
	cRightMotor = RightMotor.eMotor; //�⡼���β�ž���μ����Τ���
 	cLeftMotor = LeftMotor.eMotor; //�⡼���β�ž���μ����Τ���

};

cell tCyclicTask GetLogTask{
	cBody = GetLogTaskBody.eBody;
	cyclicAttribute = C_EXP("TA_NULL");
	cyclicTime = 20;
	cyclicPhase = 1;
	priority = 6;
	stackSize = 1024;
};

